module qnigma_tcp
  import
    qnigma_pkg::*;
(
  input  logic                  clk,
  input  logic                  rst,
  input  logic                  tick_ms,
  input  logic                  tick_s,

  input logic                   rtr_det,
  input logic                   pfx_avl,
  input logic                   dns_avl,
  input logic [15:0]            mtu,
  
  input  meta_mac_t             rx_meta_mac,
  input  meta_ip_t              rx_meta_ip,
  input  meta_tcp_t             rx_meta_tcp,
  input  meta_tcp_pres_t        rx_meta_tcp_pres,
  input  logic                  rcv,
  output meta_mac_t             tx_meta_mac,
  output meta_ip_t              tx_meta_ip,
  output meta_tcp_t             tx_meta_tcp,
  output meta_tcp_pres_t        tx_meta_tcp_pres,
  output logic                  tx_pend,
  input  logic                  tx_acpt,
  input  logic                  tx_done,
  input  logic [7:0]            dat_in,
  input  logic                  val_in,
  output logic                  cts_in,
  input  logic                  frc_in,
  output logic [7:0]            dat_out,
  output logic                  val_out,
  input  logic                  pld_req_tx,
  output logic                  pld_val_tx,
  output logic [7:0]            pld_dat_tx,
  input  logic                  pld_sof_rx,
  input  logic                  pld_val_rx,
  input  logic [7:0]            pld_dat_rx,
  input  logic                  connect_name,
  input  logic                  connect_addr,
  input  logic                  listen,
  input  logic                  disconnect,
  input  ip_t                   rem_ip,
  input  logic  [15:0]          rem_port,
  input  logic  [15:0]          loc_port,
  output logic [15:0]           con_port,
  output ip_t                   con_ip,
  output logic                  icmp_ns_req,
  input  logic                  icmp_ns_err,
  input  logic                  icmp_ns_acc,
  output ip_t                   icmp_ip_req,
  input  mac_t                  icmp_mac_rsp,
  input  logic                  icmp_rsp_ok,
  output logic                  dns_host_req,
  input  logic                  dns_host_acc,
  input  ip_t                   dns_host_addr,
  input  logic                  dns_val,
  input  logic                  dns_err,
  output tcp_stat_t             status

);

  tcp_pld_info_t tx_pld_info;

  logic send_pld;
  logic req;
  logic tcp_rst;
  logic send_ka;
  logic ka_sent;
  logic ka_dcn;
  logic flush_rx;
  logic flushed_rx;
  logic flush_tx;
  logic flushed_tx;
 
  tcp_opt_sack_t loc_sack;
  logic          send_ack;
  logic          ack_sent;

  meta_mac_t      tx_meta_mac_eng;
  meta_ip_t       tx_meta_ip_eng;
  meta_tcp_t      tx_meta_tcp_eng;
  meta_tcp_pres_t tx_meta_tcp_pres_eng;

  logic          ini;

  logic [31:0]    loc_ack;

  logic           dup_det;
  logic [31:0]    dup_ack;
  logic           soft_rst;
  logic           force_dcn;
  logic pld_sent;
  logic acpt_eng;
   
  tcb_t tcb;
  assign status = tcb.status;

  meta_mac_t meta_mac_eng;
  meta_ip_t  meta_ip_eng;
  meta_tcp_t meta_tcp_eng;
  logic      tx_pend_eng;
  /*
   * This is the global reset for all TCP-related logic
   * generated by engine based on TCP state
   */
  logic      logic_rst;
  logic flt_src_port;
  logic flt_dst_port;
  logic [31:0] last_seq;

  assign flt_src_port = rem_port == rx_meta_tcp.src;
  assign flt_dst_port = loc_port == rx_meta_tcp.dst;


  qnigma_tcp_engine qnigma_tcp_engine_inst (
    .clk              (clk                  ),
    .rst              (rst                  ),
    .logic_rst        (logic_rst            ),
    .tick_ms          (tick_ms              ),
    .rtr_det          (rtr_det              ),
    .pfx_avl          (pfx_avl              ),
    .dns_avl          (dns_avl              ),
    .mtu              (mtu                  ),
    .tcb              (tcb                  ),
    // TCP <-> RX 
    .rx_meta_mac      (rx_meta_mac          ),
    .rx_meta_ip       (rx_meta_ip           ),
    .rx_meta_tcp      (rx_meta_tcp          ),
    .rx_meta_tcp_pres (rx_meta_tcp_pres     ),
    .rcv              (rcv                  ),
    .flt_src_port     (flt_src_port         ),
    .flt_dst_port     (flt_dst_port         ),
    // TCP <-> TX
    .tx_meta_mac      (tx_meta_mac          ),
    .tx_meta_ip       (tx_meta_ip           ),
    .tx_meta_tcp      (tx_meta_tcp          ),
    .tx_meta_tcp_pres (tx_meta_tcp_pres     ),
    .tx_pend          (tx_pend              ),
    .tx_acpt          (tx_acpt              ),
    .tx_done          (tx_done              ),
    .ini              (ini                  ),
    .val_in           (val_in               ),
    .flush            (flush_tx             ),
    .flushed          (flushed_tx           ),
    .loc_ack          (loc_ack              ),
    .loc_sack         (loc_sack             ),
    .last_seq         (last_seq             ),
    .soft_rst         (soft_rst             ),
    .force_dcn        (force_dcn            ),
    .ka_dcn           (ka_dcn               ),
    // User control
    .connect_name     (connect_name         ),
    .connect_addr     (connect_addr         ),
    .listen           (listen               ),
    .disconnect       (disconnect           ),
    .rem_ip           (rem_ip               ),
    .rem_port         (rem_port             ),
    .loc_port         (loc_port             ),
    .con_port         (con_port             ),
    .con_ip           (con_ip               ),
    // TCP <-> ICMP NS
    .icmp_ns_req      (icmp_ns_req          ),
    .icmp_ns_err      (icmp_ns_err          ),
    .icmp_ns_acc      (icmp_ns_acc          ),
    .icmp_ip_req      (icmp_ip_req          ),
    .icmp_mac_rsp     (icmp_mac_rsp         ),
    .icmp_rsp_ok      (icmp_rsp_ok          ),
    // TCP <-> DNS
    .dns_host_req     (dns_host_req         ),
    .dns_host_acc     (dns_host_acc         ),
    .dns_host_addr    (dns_host_addr        ),
    .dns_val          (dns_val              ),
    .dns_err          (dns_err              ),
    
    .send_ka          (send_ka              ),
    .ka_sent          (ka_sent              ),
    .send_pld         (send_pld             ),
    .pld_info         (tx_pld_info          ),
    .pld_sent         (pld_sent             ),
    .send_ack         (send_ack             ),
    .ack_sent         (ack_sent             )
  );
  ////////////////////////////////
  // Receive buffer and control //
  ////////////////////////////////
  qnigma_tcp_rx_ctl qnigma_tcp_rx_ctl_inst (
    .clk              (clk                  ),
    .tick_ms          (tick_ms              ),
    .rst              (logic_rst            ),
    .tcb              (tcb                  ),
    .meta_tcp         (rx_meta_tcp          ),
    .rcv              (rcv                  ),
    .pld_dat          (pld_dat_rx           ),
    .pld_val          (pld_val_rx           ),
    .pld_sof          (pld_sof_rx           ),
    .dat_out          (dat_out              ),
    .val_out          (val_out              ),
    .ini              (ini                  ),
    .flush            (flush_rx             ),
    .flushed          (flushed_rx           ),
    .loc_ack          (loc_ack              ),
    .loc_sack         (loc_sack             ),
    .send_ack         (send_ack             ),
    .ack_sent         (ack_sent             )
  );

  qnigma_tcp_tx_ctl  qnigma_tcp_tx_ctl_inst (
    .clk              (clk                  ),
    .rst              (logic_rst            ),
    .dat              (dat_in               ),
    .val              (val_in               ),
    .cts              (cts_in               ),
    .frc              (frc_in               ),
    .flush            (flush_tx             ),
    .flushed          (flushed_tx           ),
    .tcb              (tcb                  ),
    .pld_val          (pld_val_tx           ),
    .pld_dat          (pld_dat_tx           ),
    .pld_req          (pld_req_tx           ),
    .ini              (ini                  ),
    .dup_ack          (dup_ack              ),
    .dup_det          (dup_det              ),
    .soft_rst         (soft_rst             ),
    .pld_info         (tx_pld_info          ),
    .send             (send_pld             ),
    .sent             (pld_sent             ),
    .force_dcn        (force_dcn            )
  );

  qnigma_tcp_ka qnigma_tcp_ka_inst (
    .clk              (clk                  ),
    .tick_s           (tick_s               ),
    .rst              (logic_rst            ),
    .tcb              (tcb                  ),
    .flt_src_port     (flt_src_port         ),
    .flt_dst_port     (flt_dst_port         ),
    .rcv              (rcv                  ),
    .send             (send_ka              ), // Send send event
    .sent             (ka_sent              ),
    .dcn              (ka_dcn               )  // Force disconnect (due to send timeout)
  );

  qnigma_tcp_fast_rtx qnigma_tcp_fast_rtx_inst (
    .clk               (clk                 ),
    .rst               (logic_rst           ),
    .tcb               (tcb                 ),
    .meta              (rx_meta_tcp         ),
    .val               (rcv                 ),
    .dup_det           (dup_det             ),
    .dup_ack           (dup_ack             ),
    .last_seq          (last_seq            )
  );

endmodule : qnigma_tcp
