module math_chacha20_poly1305_qnigma #(
  parameter int ROUNDS = 20  
) 
(
  // input  logic clk,
  // input  logic rst,
  // input  logic vi , 
  // output logic vo , // Done
  // input  cha_ada_t ada, // Associated data
  // input  cha_non_t non, // Nonce
  // input  cha_key_t key, // Key
  // output cha_tag_t tag  // Authentication tag
);

  // math_poly1305_keygen keygen_inst (
  //   .clk (clk),
  //   .rst (rst),
  //   .key (),
  //   .non (),
  //   .otk ()  // One-time key
  // );

  // qnigma_math_chacha20 chacha20_inst (
  //   .clk (clk),
  //   .rst (rst),
  //   .key (),
  //   .non ()
  // );

  // math_poly1305_mac mac_inst (
  //   .clk (clk),
  //   .rst (rst),
  //   .ada (),
  //   .otk (),
  //   .ctx ()
  // );

endmodule
