// Network top-level simulation 
module top (
  input  logic               clk                     ,
  input  logic               rst                     ,
  input  logic               phy_rx_clk              ,
  input  logic               phy_rx_err              ,
  input  logic               phy_rx_val              ,
  input  logic       [7:0]   phy_rx_dat              ,  
  output logic               phy_tx_clk              ,
  output logic               phy_tx_err              ,
  output logic               phy_tx_val              ,
  output logic       [7:0]   phy_tx_dat              ,

  input  logic       [7:0]   tcp_dat_in              ,
  input  logic               tcp_val_in              ,
  output logic               tcp_cts_in              ,
  input  logic               tcp_frc_in              ,
  output logic       [7:0]   tcp_dat_out             ,
  output logic               tcp_val_out             ,
  input  logic       [127:0] tcp_rem_ip              ,
  input  logic       [15:0]  tcp_rem_port            ,
  input  logic       [15:0]  tcp_loc_port            ,
  
  input  logic       [255:0] tcp_hostname_str        ,
  input  logic       [7:0]   tcp_hostname_len        ,
  input  logic               tcp_connect_name        ,
  input  logic               tcp_connect_addr        ,
  input  logic               tcp_listen              ,
  input  logic               tcp_disconnect          ,
  output logic       [127:0] tcp_con_ip              ,
  output logic       [15:0]  tcp_con_port            ,
 
  output logic               tcp_status_idle         ,
  output logic               tcp_status_wait_dns     ,
  output logic               tcp_status_listening    ,
  output logic               tcp_status_connecting   ,
  output logic               tcp_status_connected    ,
  output logic               tcp_status_disconnecting,
  input  logic  [15:0]       udp_len                 ,
  input  logic  [7:0]        udp_din                 ,
  input  logic               udp_vin                 ,
  output logic               udp_cts                 ,
  output logic  [7:0]        udp_dout                ,
  output logic               udp_vout                ,
  input  logic  [15:0]       udp_loc_port            ,
  output logic  [127:0]      udp_ip_rx               ,
  output logic  [15:0]       udp_rem_port_rx         ,
  input  logic  [127:0]      udp_ip_tx               ,
  input  logic  [15:0]       udp_rem_port
);

  wrap wrap (
    .clk                      (clk                      ),
    .rst                      (rst                      ),
    .phy_rx_clk               (phy_rx_clk               ),
    .phy_rx_err               (phy_rx_err               ),
    .phy_rx_val               (phy_rx_val               ),
    .phy_rx_dat               (phy_rx_dat               ),  
    .phy_tx_clk               (phy_tx_clk               ),
    .phy_tx_err               (phy_tx_err               ),
    .phy_tx_val               (phy_tx_val               ),
    .phy_tx_dat               (phy_tx_dat               ),
    .tcp_dat_in               (tcp_dat_in               ),
    .tcp_val_in               (tcp_val_in               ),
    .tcp_cts_in               (tcp_cts_in               ),
    .tcp_frc_in               (tcp_frc_in               ),
    .tcp_dat_out              (tcp_dat_out              ),
    .tcp_val_out              (tcp_val_out              ),
    .tcp_rem_ip               (tcp_rem_ip               ),
    .tcp_rem_port             (tcp_rem_port             ),
    .tcp_loc_port             (tcp_loc_port             ),
    .tcp_hostname_str         (tcp_hostname_str         ),
    .tcp_hostname_len         (tcp_hostname_len         ),
    .tcp_connect_name         (tcp_connect_name         ),
    .tcp_connect_addr         (tcp_connect_addr         ),
    .tcp_listen               (tcp_listen               ),
    .tcp_disconnect           (tcp_disconnect           ),
    .tcp_con_ip               (tcp_con_ip               ),
    .tcp_con_port             (tcp_con_port             ),
    .tcp_status_idle          (tcp_status_idle          ),
    .tcp_status_wait_dns      (tcp_status_wait_dns      ),
    .tcp_status_listening     (tcp_status_listening     ),
    .tcp_status_connecting    (tcp_status_connecting    ),
    .tcp_status_connected     (tcp_status_connected     ),
    .tcp_status_disconnecting (tcp_status_disconnecting ),
    .udp_len                  (udp_len                  ),
    .udp_din                  (udp_din                  ),
    .udp_vin                  (udp_vin                  ),
    .udp_cts                  (udp_cts                  ),
    .udp_dout                 (udp_dout                 ),
    .udp_vout                 (udp_vout                 ),
    .udp_loc_port             (udp_loc_port             ),
    .udp_ip_rx                (udp_ip_rx                ),
    .udp_rem_port_rx          (udp_rem_port_rx          ),
    .udp_ip_tx                (udp_ip_tx                ),
    .udp_rem_port             (udp_rem_port             )
  );

endmodule : top
