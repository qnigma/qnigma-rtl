localparam REFCLK_HZ = 12500;